�� sr proiect.logic.GameStatel�K���� I bugetL coadat Ljava/util/Queue;L hotelt Lproiect/model/Hotel;xp ��sr java.util.LinkedList)S]J`�"  xpw    xsr proiect.model.Hotel[`�~��d L cameret Ljava/util/Set;xpsr java.util.LinkedHashSet�l�Z��*  xr java.util.HashSet�D�����4  xpw   ?@     sr proiect.model.CameraW�JO\�/ L clientt Lproiect/model/Client;L tipt Lproiect/model/TipCamera;xpsr proiect.model.Client_��뫊� I 	nrAnimaleI nrDaysL numet Ljava/lang/String;xp      t Ghita~r proiect.model.TipCamera          xr java.lang.Enum          xpt DOUBLEsq ~ sq ~       q ~ q ~ sq ~ sq ~       q ~ q ~ sq ~ sq ~       q ~ q ~ sq ~ sq ~       t Ghitaq ~ sq ~ sq ~       q ~  q ~ sq ~ pq ~ sq ~ sq ~       q ~  q ~ x