�� sr proiect.logic.GameStatel�K���� L bugett +Ljava/util/concurrent/atomic/AtomicInteger;L coadat Ljava/util/Queue;L hotelt Lproiect/model/Hotel;xpsr )java.util.concurrent.atomic.AtomicIntegerV?^̌l� I valuexr java.lang.Number������  xp B@sr java.util.LinkedList)S]J`�"  xpw   sr proiect.model.Client_��뫊� I 	nrAnimaleI nrDaysL numet Ljava/lang/String;xp      t Ghitasq ~ 
      q ~ sq ~ 
      q ~ xsr proiect.model.Hotel[`�~��d L cameret Ljava/util/Set;xpsr java.util.LinkedHashSet�l�Z��*  xr java.util.HashSet�D�����4  xpw   ?@      x